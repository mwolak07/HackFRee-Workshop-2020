
//
// Verific Verilog Description of module top_module
//

module top_module (pll_LOCKED, pll_CLK, btn1, led1, led2);
    input pll_LOCKED /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input pll_CLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input btn1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output led1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output led2 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    
    wire n487 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n555 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n519 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n515 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n587 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n551 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n511 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n507 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n583 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n547 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n503 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n499 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n579 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n543 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n495 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n491 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n575 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n539 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n571 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n535 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n567 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n531 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n563 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n527 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n559 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    wire n523 /* verific EFX_ATTRIBUTE__IS_CMB_LOOP_NET=TRUE */ ;
    
    wire n207, n218, n229, n240, n251, n262, n273, n284, n295, 
        n306, n317, n328, n339, n350, n361, n372, n383, n394, 
        n405, n416, n427, n438, n449, n460, n471, n482, n33, 
        n34, n36, n40, n41, n43, n47, n48, n50, n54, n55, 
        n57, n60, n61, n62, n63, n64, n65, n66, n67, n70, 
        n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, 
        n81, n82, n83, n84, n87, n88, n89, n90, n91, n92, 
        n93, n94, n95, n96, n97, n98, n99, n100, n101, n104, 
        n105, n106, n107, n108, n109, n110, n111, n112, n113, 
        n114, n115, n116, n117, n118, n121, n122, n123, n124, 
        n125, n126, n127, n128, n129, n130, n189, n190, n191, 
        n192, n194, n195, n199, n200, n201, n202, n204, n205, 
        n209, n210, n211, n212, n214, n215, n219, n220, n221, 
        n222, n224, n225, n228, n229_2, n232, n233, n238, n239, 
        n246, n247, n252, n253, n258, n259, n266, n267, n272, 
        n273_2, n278, n279, n286, n287, n292, n293, n298, n299, 
        n306_2, n307, \pll_CLK~O , n312, n313;
    
    EFX_FF \n207~FF  (.D(n33), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n207~FF .CLK_POLARITY = 1'b1;
    defparam \n207~FF .CE_POLARITY = 1'b1;
    defparam \n207~FF .SR_POLARITY = 1'b0;
    defparam \n207~FF .D_POLARITY = 1'b1;
    defparam \n207~FF .SR_SYNC = 1'b0;
    defparam \n207~FF .SR_VALUE = 1'b0;
    defparam \n207~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n218~FF  (.D(n34), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n218~FF .CLK_POLARITY = 1'b1;
    defparam \n218~FF .CE_POLARITY = 1'b1;
    defparam \n218~FF .SR_POLARITY = 1'b0;
    defparam \n218~FF .D_POLARITY = 1'b1;
    defparam \n218~FF .SR_SYNC = 1'b0;
    defparam \n218~FF .SR_VALUE = 1'b0;
    defparam \n218~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n229~FF  (.D(n36), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n229~FF .CLK_POLARITY = 1'b1;
    defparam \n229~FF .CE_POLARITY = 1'b1;
    defparam \n229~FF .SR_POLARITY = 1'b0;
    defparam \n229~FF .D_POLARITY = 1'b1;
    defparam \n229~FF .SR_SYNC = 1'b0;
    defparam \n229~FF .SR_VALUE = 1'b0;
    defparam \n229~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n240~FF  (.D(n40), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n240~FF .CLK_POLARITY = 1'b1;
    defparam \n240~FF .CE_POLARITY = 1'b1;
    defparam \n240~FF .SR_POLARITY = 1'b0;
    defparam \n240~FF .D_POLARITY = 1'b1;
    defparam \n240~FF .SR_SYNC = 1'b0;
    defparam \n240~FF .SR_VALUE = 1'b0;
    defparam \n240~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n251~FF  (.D(n41), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n251~FF .CLK_POLARITY = 1'b1;
    defparam \n251~FF .CE_POLARITY = 1'b1;
    defparam \n251~FF .SR_POLARITY = 1'b0;
    defparam \n251~FF .D_POLARITY = 1'b1;
    defparam \n251~FF .SR_SYNC = 1'b0;
    defparam \n251~FF .SR_VALUE = 1'b0;
    defparam \n251~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n262~FF  (.D(n43), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n262~FF .CLK_POLARITY = 1'b1;
    defparam \n262~FF .CE_POLARITY = 1'b1;
    defparam \n262~FF .SR_POLARITY = 1'b0;
    defparam \n262~FF .D_POLARITY = 1'b1;
    defparam \n262~FF .SR_SYNC = 1'b0;
    defparam \n262~FF .SR_VALUE = 1'b0;
    defparam \n262~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n273~FF  (.D(n47), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n273~FF .CLK_POLARITY = 1'b1;
    defparam \n273~FF .CE_POLARITY = 1'b1;
    defparam \n273~FF .SR_POLARITY = 1'b0;
    defparam \n273~FF .D_POLARITY = 1'b1;
    defparam \n273~FF .SR_SYNC = 1'b0;
    defparam \n273~FF .SR_VALUE = 1'b0;
    defparam \n273~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n284~FF  (.D(n48), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n284~FF .CLK_POLARITY = 1'b1;
    defparam \n284~FF .CE_POLARITY = 1'b1;
    defparam \n284~FF .SR_POLARITY = 1'b0;
    defparam \n284~FF .D_POLARITY = 1'b1;
    defparam \n284~FF .SR_SYNC = 1'b0;
    defparam \n284~FF .SR_VALUE = 1'b0;
    defparam \n284~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n295~FF  (.D(n50), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n295~FF .CLK_POLARITY = 1'b1;
    defparam \n295~FF .CE_POLARITY = 1'b1;
    defparam \n295~FF .SR_POLARITY = 1'b0;
    defparam \n295~FF .D_POLARITY = 1'b1;
    defparam \n295~FF .SR_SYNC = 1'b0;
    defparam \n295~FF .SR_VALUE = 1'b0;
    defparam \n295~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n306~FF  (.D(n54), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n306~FF .CLK_POLARITY = 1'b1;
    defparam \n306~FF .CE_POLARITY = 1'b1;
    defparam \n306~FF .SR_POLARITY = 1'b0;
    defparam \n306~FF .D_POLARITY = 1'b1;
    defparam \n306~FF .SR_SYNC = 1'b0;
    defparam \n306~FF .SR_VALUE = 1'b0;
    defparam \n306~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n317~FF  (.D(n55), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n317~FF .CLK_POLARITY = 1'b1;
    defparam \n317~FF .CE_POLARITY = 1'b1;
    defparam \n317~FF .SR_POLARITY = 1'b0;
    defparam \n317~FF .D_POLARITY = 1'b1;
    defparam \n317~FF .SR_SYNC = 1'b0;
    defparam \n317~FF .SR_VALUE = 1'b0;
    defparam \n317~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n328~FF  (.D(n57), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n328~FF .CLK_POLARITY = 1'b1;
    defparam \n328~FF .CE_POLARITY = 1'b1;
    defparam \n328~FF .SR_POLARITY = 1'b0;
    defparam \n328~FF .D_POLARITY = 1'b1;
    defparam \n328~FF .SR_SYNC = 1'b0;
    defparam \n328~FF .SR_VALUE = 1'b0;
    defparam \n328~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n339~FF  (.D(n60), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n339~FF .CLK_POLARITY = 1'b1;
    defparam \n339~FF .CE_POLARITY = 1'b1;
    defparam \n339~FF .SR_POLARITY = 1'b0;
    defparam \n339~FF .D_POLARITY = 1'b1;
    defparam \n339~FF .SR_SYNC = 1'b0;
    defparam \n339~FF .SR_VALUE = 1'b0;
    defparam \n339~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n350~FF  (.D(n62), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n350~FF .CLK_POLARITY = 1'b1;
    defparam \n350~FF .CE_POLARITY = 1'b1;
    defparam \n350~FF .SR_POLARITY = 1'b0;
    defparam \n350~FF .D_POLARITY = 1'b1;
    defparam \n350~FF .SR_SYNC = 1'b0;
    defparam \n350~FF .SR_VALUE = 1'b0;
    defparam \n350~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n361~FF  (.D(n67), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n361~FF .CLK_POLARITY = 1'b1;
    defparam \n361~FF .CE_POLARITY = 1'b1;
    defparam \n361~FF .SR_POLARITY = 1'b0;
    defparam \n361~FF .D_POLARITY = 1'b1;
    defparam \n361~FF .SR_SYNC = 1'b0;
    defparam \n361~FF .SR_VALUE = 1'b0;
    defparam \n361~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n372~FF  (.D(n74), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n372~FF .CLK_POLARITY = 1'b1;
    defparam \n372~FF .CE_POLARITY = 1'b1;
    defparam \n372~FF .SR_POLARITY = 1'b0;
    defparam \n372~FF .D_POLARITY = 1'b1;
    defparam \n372~FF .SR_SYNC = 1'b0;
    defparam \n372~FF .SR_VALUE = 1'b0;
    defparam \n372~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n383~FF  (.D(n79), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n383~FF .CLK_POLARITY = 1'b1;
    defparam \n383~FF .CE_POLARITY = 1'b1;
    defparam \n383~FF .SR_POLARITY = 1'b0;
    defparam \n383~FF .D_POLARITY = 1'b1;
    defparam \n383~FF .SR_SYNC = 1'b0;
    defparam \n383~FF .SR_VALUE = 1'b0;
    defparam \n383~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n394~FF  (.D(n84), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n394~FF .CLK_POLARITY = 1'b1;
    defparam \n394~FF .CE_POLARITY = 1'b1;
    defparam \n394~FF .SR_POLARITY = 1'b0;
    defparam \n394~FF .D_POLARITY = 1'b1;
    defparam \n394~FF .SR_SYNC = 1'b0;
    defparam \n394~FF .SR_VALUE = 1'b0;
    defparam \n394~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n405~FF  (.D(n91), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n405~FF .CLK_POLARITY = 1'b1;
    defparam \n405~FF .CE_POLARITY = 1'b1;
    defparam \n405~FF .SR_POLARITY = 1'b0;
    defparam \n405~FF .D_POLARITY = 1'b1;
    defparam \n405~FF .SR_SYNC = 1'b0;
    defparam \n405~FF .SR_VALUE = 1'b0;
    defparam \n405~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n416~FF  (.D(n96), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n416~FF .CLK_POLARITY = 1'b1;
    defparam \n416~FF .CE_POLARITY = 1'b1;
    defparam \n416~FF .SR_POLARITY = 1'b0;
    defparam \n416~FF .D_POLARITY = 1'b1;
    defparam \n416~FF .SR_SYNC = 1'b0;
    defparam \n416~FF .SR_VALUE = 1'b0;
    defparam \n416~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n427~FF  (.D(n101), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n427~FF .CLK_POLARITY = 1'b1;
    defparam \n427~FF .CE_POLARITY = 1'b1;
    defparam \n427~FF .SR_POLARITY = 1'b0;
    defparam \n427~FF .D_POLARITY = 1'b1;
    defparam \n427~FF .SR_SYNC = 1'b0;
    defparam \n427~FF .SR_VALUE = 1'b0;
    defparam \n427~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n438~FF  (.D(n108), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n438~FF .CLK_POLARITY = 1'b1;
    defparam \n438~FF .CE_POLARITY = 1'b1;
    defparam \n438~FF .SR_POLARITY = 1'b0;
    defparam \n438~FF .D_POLARITY = 1'b1;
    defparam \n438~FF .SR_SYNC = 1'b0;
    defparam \n438~FF .SR_VALUE = 1'b0;
    defparam \n438~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n449~FF  (.D(n113), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n449~FF .CLK_POLARITY = 1'b1;
    defparam \n449~FF .CE_POLARITY = 1'b1;
    defparam \n449~FF .SR_POLARITY = 1'b0;
    defparam \n449~FF .D_POLARITY = 1'b1;
    defparam \n449~FF .SR_SYNC = 1'b0;
    defparam \n449~FF .SR_VALUE = 1'b0;
    defparam \n449~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n460~FF  (.D(n118), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n460~FF .CLK_POLARITY = 1'b1;
    defparam \n460~FF .CE_POLARITY = 1'b1;
    defparam \n460~FF .SR_POLARITY = 1'b0;
    defparam \n460~FF .D_POLARITY = 1'b1;
    defparam \n460~FF .SR_SYNC = 1'b0;
    defparam \n460~FF .SR_VALUE = 1'b0;
    defparam \n460~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n471~FF  (.D(n125), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n471~FF .CLK_POLARITY = 1'b1;
    defparam \n471~FF .CE_POLARITY = 1'b1;
    defparam \n471~FF .SR_POLARITY = 1'b0;
    defparam \n471~FF .D_POLARITY = 1'b1;
    defparam \n471~FF .SR_SYNC = 1'b0;
    defparam \n471~FF .SR_VALUE = 1'b0;
    defparam \n471~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \n482~FF  (.D(n130), .CE(1'b1), .CLK(\pll_CLK~O ), .SR(btn1), 
           .Q(n482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(14)
    defparam \n482~FF .CLK_POLARITY = 1'b1;
    defparam \n482~FF .CE_POLARITY = 1'b1;
    defparam \n482~FF .SR_POLARITY = 1'b0;
    defparam \n482~FF .D_POLARITY = 1'b1;
    defparam \n482~FF .SR_SYNC = 1'b0;
    defparam \n482~FF .SR_VALUE = 1'b0;
    defparam \n482~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 i120 (.I1(n36), .I2(n194), .I3(n195), .O(n36)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i120.LUTMASK = 16'h00FC;
    EFX_LUT4 i130 (.I1(n40), .I2(n199), .I3(n200), .O(n40)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i130.LUTMASK = 16'h00FC;
    EFX_LUT4 i140 (.I1(n41), .I2(n201), .I3(n202), .O(n41)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i140.LUTMASK = 16'h00FC;
    EFX_LUT4 i150 (.I1(n43), .I2(n204), .I3(n205), .O(n43)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i150.LUTMASK = 16'h00FC;
    EFX_LUT4 i160 (.I1(n47), .I2(n209), .I3(n210), .O(n47)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i160.LUTMASK = 16'h00FC;
    EFX_LUT4 i170 (.I1(n48), .I2(n211), .I3(n212), .O(n48)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i170.LUTMASK = 16'h00FC;
    EFX_LUT4 i180 (.I1(n50), .I2(n214), .I3(n215), .O(n50)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i180.LUTMASK = 16'h00FC;
    EFX_LUT4 i190 (.I1(n54), .I2(n219), .I3(n220), .O(n54)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i190.LUTMASK = 16'h00FC;
    EFX_LUT4 i200 (.I1(n55), .I2(n221), .I3(n222), .O(n55)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i200.LUTMASK = 16'h00FC;
    EFX_LUT4 i210 (.I1(n57), .I2(n224), .I3(n225), .O(n57)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i210.LUTMASK = 16'h00FC;
    EFX_LUT4 i220 (.I1(n60), .I2(n228), .I3(n229_2), .O(n60)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i220.LUTMASK = 16'h00FC;
    EFX_LUT4 i230 (.I1(n62), .I2(n232), .I3(n233), .O(n62)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i230.LUTMASK = 16'h00FC;
    EFX_LUT4 i240 (.I1(n67), .I2(n238), .I3(n239), .O(n67)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i240.LUTMASK = 16'h00FC;
    EFX_LUT4 i250 (.I1(n74), .I2(n246), .I3(n247), .O(n74)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i250.LUTMASK = 16'h00FC;
    EFX_LUT4 i260 (.I1(n79), .I2(n252), .I3(n253), .O(n79)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i260.LUTMASK = 16'h00FC;
    EFX_LUT4 i270 (.I1(n84), .I2(n258), .I3(n259), .O(n84)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i270.LUTMASK = 16'h00FC;
    EFX_LUT4 i280 (.I1(n91), .I2(n266), .I3(n267), .O(n91)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i280.LUTMASK = 16'h00FC;
    EFX_LUT4 i290 (.I1(n96), .I2(n272), .I3(n273_2), .O(n96)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i290.LUTMASK = 16'h00FC;
    EFX_LUT4 i300 (.I1(n101), .I2(n278), .I3(n279), .O(n101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i300.LUTMASK = 16'h00FC;
    EFX_LUT4 i310 (.I1(n108), .I2(n286), .I3(n287), .O(n108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i310.LUTMASK = 16'h00FC;
    EFX_LUT4 i320 (.I1(n113), .I2(n292), .I3(n293), .O(n113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i320.LUTMASK = 16'h00FC;
    EFX_LUT4 i330 (.I1(n118), .I2(n298), .I3(n299), .O(n118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i330.LUTMASK = 16'h00FC;
    EFX_LUT4 i340 (.I1(n125), .I2(n306_2), .I3(n307), .O(n125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i340.LUTMASK = 16'h00FC;
    EFX_LUT4 i350 (.I1(n130), .I2(n312), .I3(n313), .O(n130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i350.LUTMASK = 16'h00FC;
    EFX_LUT4 LUT__446 (.I0(n487), .I1(n491), .O(led1)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__446.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__447 (.I0(n61), .I1(n487), .I2(btn1), .I3(pll_LOCKED), 
            .O(n313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__447.LUTMASK = 16'h0503;
    EFX_ADD \add_8/i26  (.I0(n487), .I1(1'b0), .CI(n64), .O(n61)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i26 .I0_POLARITY = 1'b1;
    defparam \add_8/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i25  (.I0(n491), .I1(1'b0), .CI(n66), .O(n63), .CO(n64)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i25 .I0_POLARITY = 1'b1;
    defparam \add_8/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i24  (.I0(n495), .I1(1'b0), .CI(n71), .O(n65), .CO(n66)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i24 .I0_POLARITY = 1'b1;
    defparam \add_8/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i23  (.I0(n499), .I1(1'b0), .CI(n73), .O(n70), .CO(n71)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i23 .I0_POLARITY = 1'b1;
    defparam \add_8/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i22  (.I0(n503), .I1(1'b0), .CI(n76), .O(n72), .CO(n73)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i22 .I0_POLARITY = 1'b1;
    defparam \add_8/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i21  (.I0(n507), .I1(1'b0), .CI(n78), .O(n75), .CO(n76)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i21 .I0_POLARITY = 1'b1;
    defparam \add_8/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i20  (.I0(n511), .I1(1'b0), .CI(n81), .O(n77), .CO(n78)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i20 .I0_POLARITY = 1'b1;
    defparam \add_8/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i19  (.I0(n515), .I1(1'b0), .CI(n83), .O(n80), .CO(n81)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i19 .I0_POLARITY = 1'b1;
    defparam \add_8/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i18  (.I0(n519), .I1(1'b0), .CI(n88), .O(n82), .CO(n83)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i18 .I0_POLARITY = 1'b1;
    defparam \add_8/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i17  (.I0(n523), .I1(1'b0), .CI(n90), .O(n87), .CO(n88)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i17 .I0_POLARITY = 1'b1;
    defparam \add_8/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i16  (.I0(n527), .I1(1'b0), .CI(n93), .O(n89), .CO(n90)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i16 .I0_POLARITY = 1'b1;
    defparam \add_8/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i15  (.I0(n531), .I1(1'b0), .CI(n95), .O(n92), .CO(n93)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i15 .I0_POLARITY = 1'b1;
    defparam \add_8/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i14  (.I0(n535), .I1(1'b0), .CI(n98), .O(n94), .CO(n95)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i14 .I0_POLARITY = 1'b1;
    defparam \add_8/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i13  (.I0(n539), .I1(1'b0), .CI(n100), .O(n97), .CO(n98)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i13 .I0_POLARITY = 1'b1;
    defparam \add_8/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i12  (.I0(n543), .I1(1'b0), .CI(n105), .O(n99), .CO(n100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i12 .I0_POLARITY = 1'b1;
    defparam \add_8/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i11  (.I0(n547), .I1(1'b0), .CI(n107), .O(n104), 
            .CO(n105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i11 .I0_POLARITY = 1'b1;
    defparam \add_8/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i10  (.I0(n551), .I1(1'b0), .CI(n110), .O(n106), 
            .CO(n107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i10 .I0_POLARITY = 1'b1;
    defparam \add_8/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i9  (.I0(n555), .I1(1'b0), .CI(n112), .O(n109), .CO(n110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i9 .I0_POLARITY = 1'b1;
    defparam \add_8/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i8  (.I0(n559), .I1(1'b0), .CI(n115), .O(n111), .CO(n112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i8 .I0_POLARITY = 1'b1;
    defparam \add_8/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i7  (.I0(n563), .I1(1'b0), .CI(n117), .O(n114), .CO(n115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i7 .I0_POLARITY = 1'b1;
    defparam \add_8/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i6  (.I0(n567), .I1(1'b0), .CI(n122), .O(n116), .CO(n117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i6 .I0_POLARITY = 1'b1;
    defparam \add_8/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i5  (.I0(n571), .I1(1'b0), .CI(n124), .O(n121), .CO(n122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i5 .I0_POLARITY = 1'b1;
    defparam \add_8/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i4  (.I0(n575), .I1(1'b0), .CI(n127), .O(n123), .CO(n124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i4 .I0_POLARITY = 1'b1;
    defparam \add_8/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i3  (.I0(n579), .I1(1'b0), .CI(n129), .O(n126), .CO(n127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i3 .I0_POLARITY = 1'b1;
    defparam \add_8/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \add_8/i2  (.I0(n583), .I1(n587), .CI(1'b0), .O(n128), .CO(n129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/mwola/OneDrive/Coding/2020/HackFRee-Workshop-2020/PllClkExample/top.v(13)
    defparam \add_8/i2 .I0_POLARITY = 1'b1;
    defparam \add_8/i2 .I1_POLARITY = 1'b1;
    EFX_LUT4 LUT__448 (.I0(n61), .I1(n487), .I2(btn1), .I3(pll_LOCKED), 
            .O(n312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__448.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__449 (.I0(btn1), .I1(n482), .I2(n130), .I3(n313), .O(n487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__449.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__450 (.I0(n109), .I1(n555), .I2(btn1), .I3(pll_LOCKED), 
            .O(n215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__450.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__451 (.I0(n109), .I1(n555), .I2(btn1), .I3(pll_LOCKED), 
            .O(n214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__451.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__452 (.I0(btn1), .I1(n295), .I2(n50), .I3(n215), .O(n555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__452.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__453 (.I0(n82), .I1(n519), .I2(btn1), .I3(pll_LOCKED), 
            .O(n259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__453.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__454 (.I0(n82), .I1(n519), .I2(btn1), .I3(pll_LOCKED), 
            .O(n258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__454.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__455 (.I0(btn1), .I1(n394), .I2(n84), .I3(n259), .O(n519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__455.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__456 (.I0(btn1), .I1(pll_LOCKED), .I2(n587), .O(n189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__456.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__457 (.I0(btn1), .I1(pll_LOCKED), .I2(n587), .O(n190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141 */ ;
    defparam LUT__457.LUTMASK = 16'h4141;
    EFX_LUT4 LUT__458 (.I0(n128), .I1(n583), .I2(btn1), .I3(pll_LOCKED), 
            .O(n191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__458.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__459 (.I0(n128), .I1(n583), .I2(btn1), .I3(pll_LOCKED), 
            .O(n192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__459.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__460 (.I0(n80), .I1(n515), .I2(btn1), .I3(pll_LOCKED), 
            .O(n267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__460.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__461 (.I0(n80), .I1(n515), .I2(btn1), .I3(pll_LOCKED), 
            .O(n266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__461.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__462 (.I0(btn1), .I1(n405), .I2(n91), .I3(n267), .O(n515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__462.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__463 (.I0(n126), .I1(n579), .I2(btn1), .I3(pll_LOCKED), 
            .O(n194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__463.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__464 (.I0(n126), .I1(n579), .I2(btn1), .I3(pll_LOCKED), 
            .O(n195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__464.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__465 (.I0(btn1), .I1(n207), .I2(n33), .I3(n190), .O(n587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__465.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__466 (.I0(n106), .I1(n551), .I2(btn1), .I3(pll_LOCKED), 
            .O(n220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__466.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__467 (.I0(n106), .I1(n551), .I2(btn1), .I3(pll_LOCKED), 
            .O(n219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__467.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__468 (.I0(btn1), .I1(n306), .I2(n54), .I3(n220), .O(n551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__468.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__469 (.I0(n77), .I1(n511), .I2(btn1), .I3(pll_LOCKED), 
            .O(n273_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__469.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__470 (.I0(n77), .I1(n511), .I2(btn1), .I3(pll_LOCKED), 
            .O(n272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__470.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__471 (.I0(btn1), .I1(n416), .I2(n96), .I3(n273_2), 
            .O(n511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__471.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__472 (.I0(n123), .I1(n575), .I2(btn1), .I3(pll_LOCKED), 
            .O(n199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__472.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__473 (.I0(n123), .I1(n575), .I2(btn1), .I3(pll_LOCKED), 
            .O(n200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__473.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__474 (.I0(n121), .I1(n571), .I2(btn1), .I3(pll_LOCKED), 
            .O(n201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__474.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__475 (.I0(n121), .I1(n571), .I2(btn1), .I3(pll_LOCKED), 
            .O(n202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__475.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__476 (.I0(n75), .I1(n507), .I2(btn1), .I3(pll_LOCKED), 
            .O(n279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__476.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__477 (.I0(n75), .I1(n507), .I2(btn1), .I3(pll_LOCKED), 
            .O(n278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__477.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__478 (.I0(btn1), .I1(n427), .I2(n101), .I3(n279), .O(n507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__478.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__479 (.I0(n116), .I1(n567), .I2(btn1), .I3(pll_LOCKED), 
            .O(n204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__479.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__480 (.I0(n116), .I1(n567), .I2(btn1), .I3(pll_LOCKED), 
            .O(n205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__480.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__481 (.I0(btn1), .I1(n218), .I2(n34), .I3(n192), .O(n583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__481.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__482 (.I0(n104), .I1(n547), .I2(btn1), .I3(pll_LOCKED), 
            .O(n222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__482.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__483 (.I0(n104), .I1(n547), .I2(btn1), .I3(pll_LOCKED), 
            .O(n221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__483.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__484 (.I0(btn1), .I1(n317), .I2(n55), .I3(n222), .O(n547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__484.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__485 (.I0(n72), .I1(n503), .I2(btn1), .I3(pll_LOCKED), 
            .O(n287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__485.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__486 (.I0(n72), .I1(n503), .I2(btn1), .I3(pll_LOCKED), 
            .O(n286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__486.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__487 (.I0(btn1), .I1(n438), .I2(n108), .I3(n287), .O(n503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__487.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__488 (.I0(n114), .I1(n563), .I2(btn1), .I3(pll_LOCKED), 
            .O(n209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__488.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__489 (.I0(n114), .I1(n563), .I2(btn1), .I3(pll_LOCKED), 
            .O(n210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__489.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__490 (.I0(n111), .I1(n559), .I2(btn1), .I3(pll_LOCKED), 
            .O(n211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__490.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__491 (.I0(n111), .I1(n559), .I2(btn1), .I3(pll_LOCKED), 
            .O(n212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__491.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__492 (.I0(n70), .I1(n499), .I2(btn1), .I3(pll_LOCKED), 
            .O(n293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__492.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__493 (.I0(n70), .I1(n499), .I2(btn1), .I3(pll_LOCKED), 
            .O(n292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__493.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__494 (.I0(btn1), .I1(n449), .I2(n113), .I3(n293), .O(n499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__494.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__495 (.I0(btn1), .I1(n229), .I2(n36), .I3(n195), .O(n579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__495.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__496 (.I0(n99), .I1(n543), .I2(btn1), .I3(pll_LOCKED), 
            .O(n225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__496.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__497 (.I0(n99), .I1(n543), .I2(btn1), .I3(pll_LOCKED), 
            .O(n224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__497.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__498 (.I0(btn1), .I1(n328), .I2(n57), .I3(n225), .O(n543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__498.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__499 (.I0(n65), .I1(n495), .I2(btn1), .I3(pll_LOCKED), 
            .O(n299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__499.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__500 (.I0(n65), .I1(n495), .I2(btn1), .I3(pll_LOCKED), 
            .O(n298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__500.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__501 (.I0(btn1), .I1(n460), .I2(n118), .I3(n299), .O(n495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__501.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__502 (.I0(n63), .I1(n491), .I2(btn1), .I3(pll_LOCKED), 
            .O(n307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__502.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__503 (.I0(n63), .I1(n491), .I2(btn1), .I3(pll_LOCKED), 
            .O(n306_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__503.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__504 (.I0(btn1), .I1(n471), .I2(n125), .I3(n307), .O(n491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__504.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__505 (.I0(btn1), .I1(n240), .I2(n40), .I3(n200), .O(n575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__505.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__506 (.I0(n97), .I1(n539), .I2(btn1), .I3(pll_LOCKED), 
            .O(n229_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__506.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__507 (.I0(n97), .I1(n539), .I2(btn1), .I3(pll_LOCKED), 
            .O(n228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__507.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__508 (.I0(btn1), .I1(n339), .I2(n60), .I3(n229_2), 
            .O(n539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__508.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__509 (.I0(n94), .I1(n535), .I2(btn1), .I3(pll_LOCKED), 
            .O(n232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__509.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__510 (.I0(n94), .I1(n535), .I2(btn1), .I3(pll_LOCKED), 
            .O(n233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__510.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__511 (.I0(n92), .I1(n531), .I2(btn1), .I3(pll_LOCKED), 
            .O(n238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__511.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__512 (.I0(n92), .I1(n531), .I2(btn1), .I3(pll_LOCKED), 
            .O(n239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__512.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__513 (.I0(btn1), .I1(n251), .I2(n41), .I3(n202), .O(n571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__513.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__514 (.I0(btn1), .I1(n350), .I2(n62), .I3(n233), .O(n535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__514.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__515 (.I0(n89), .I1(n527), .I2(btn1), .I3(pll_LOCKED), 
            .O(n246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__515.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__516 (.I0(n89), .I1(n527), .I2(btn1), .I3(pll_LOCKED), 
            .O(n247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__516.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__517 (.I0(n87), .I1(n523), .I2(btn1), .I3(pll_LOCKED), 
            .O(n252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__517.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__518 (.I0(n87), .I1(n523), .I2(btn1), .I3(pll_LOCKED), 
            .O(n253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__518.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__519 (.I0(btn1), .I1(n262), .I2(n43), .I3(n205), .O(n567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__519.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__520 (.I0(btn1), .I1(n361), .I2(n67), .I3(n239), .O(n531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__520.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__521 (.I0(btn1), .I1(n273), .I2(n47), .I3(n210), .O(n563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__521.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__522 (.I0(btn1), .I1(n372), .I2(n74), .I3(n247), .O(n527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__522.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__523 (.I0(btn1), .I1(n284), .I2(n48), .I3(n212), .O(n559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__523.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__524 (.I0(btn1), .I1(n383), .I2(n79), .I3(n253), .O(n523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__524.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__527 (.I0(led1), .O(led2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__527.LUTMASK = 16'h5555;
    EFX_LUT4 i100 (.I1(n33), .I2(n189), .I3(n190), .O(n33)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i100.LUTMASK = 16'h00FC;
    EFX_LUT4 i110 (.I1(n34), .I2(n191), .I3(n192), .O(n34)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i110.LUTMASK = 16'h00FC;
    EFX_GBUFCE CLKBUF__0 (.CE(1'b1), .I(pll_CLK), .O(\pll_CLK~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__0.CE_POLARITY = 1'b1;
    
endmodule

//
// Verific Verilog Description of module EFX_FF0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT410
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT411
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT412
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT413
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT414
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT415
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT416
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT417
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT418
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT419
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT420
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT421
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT422
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT423
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT424
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT425
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT426
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT427
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT428
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT429
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT430
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT431
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT432
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT433
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT434
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT435
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT436
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT437
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT438
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT439
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT440
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT441
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT442
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT443
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT444
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT445
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT446
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT447
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT448
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT449
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT450
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT451
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT452
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT453
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT454
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT455
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT456
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT457
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT458
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT459
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT460
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT461
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT462
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT463
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT464
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT465
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT466
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT467
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT468
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT469
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT470
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT471
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT472
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT473
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT474
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT475
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT476
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT477
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT478
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT479
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT480
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT481
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT482
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT483
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT484
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT485
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT486
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT487
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT488
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT489
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT490
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT491
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT492
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT493
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT494
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT495
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT496
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT497
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT498
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT499
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE0
// module not written out since it is a black box. 
//


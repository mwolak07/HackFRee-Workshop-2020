
// Efinity Top-level template
// Version: 2019.3.272
// Date: 2020-01-18 13:28

// Copyright (C) 2017 - 2019 Efinix Inc. All rights reserved.

// This file may be used as a starting point for Efinity synthesis top-level target.
// The port list here matches what is expected by Efinity constraint files generated
// by the Efinity Interface Designer.

// To use this:
//     #1)  Save this file with a different name to a different directory, where source files are kept.
//              Example: you may wish to save as C:\Users\mwola\OneDrive\Coding\2020\HackFRee-Workshop-2020\BasicExample\BasicExample.v
//     #2)  Add the newly saved file into Efinity project as design file
//     #3)  Edit the top level entity in Efinity project to:  BasicExample
//     #4)  Insert design content.


module BasicExample
(
  input clk,
  input btn1,
  input btn2,
  output led1,
  output led2
);


endmodule

